module FPGA #(
    parameter  = 
) (
    input   wire                    clk     ,
    input   wire                    rst_n   ,
    input   wire                          ,
    output  wire                          ,      
    output  reg                                 
);
//==============================================================================
// Constant Definition :
//==============================================================================




//==============================================================================
// Variable Definition :
//==============================================================================





//==============================================================================
// Logic Design :
//==============================================================================
assign 





//==============================================================================
// Sub-Module :
//==============================================================================



endmodule